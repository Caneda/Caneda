process(D, EN)
begin
   if(EN = '1') then
      Q <= D;
   end if;
end process;
