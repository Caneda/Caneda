always @ (D or EN) begin
   if (EN) begin
      Q <= D;
   end
end
