process (A, B, ...)
begin
   -- Concurrent asignments
   ...

end process;
