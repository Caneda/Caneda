always @ ( A, B, ... ) begin
   // Concurrent assignments
   ...
end
