always @ ( posedge clk ) begin
   Q <= D;
end
