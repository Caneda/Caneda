if(CONDITION) then
   -- Concurrent asignments
   ...
elsif(CONDITION) then
   -- Concurrent asignments
   ...
end if;
