signal name: TYPE;
