// name can be any name chosen for this module
module name ( A, B, X, Y, ... );

   // Constants
   parameter cons1 = VALUE;
   parameter cons2 = VALUE;
   ...

   // Inputs and outputs
   input  A, B;
   output X, Y;
   ...

   // Data types
   wire A, B;
   reg  X, Y;
   ...

   // Always statements and continous assignments
   ...

endmodule
