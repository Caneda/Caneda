-- name can be any name chosen for this architecture
-- entity is the name of the entity previously defined
ARCHITECTURE name OF entity IS
   -- Signal, component, type and constant declarations go here
   ...

BEGIN
   -- Concurrent statements and processes go here
   ...

END name;
