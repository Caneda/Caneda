-- name can be any name chosen for this package
PACKAGE name IS
   -- Constructs declaration go here
   -- Signal, component, type and constant declarations go here
   ...

END name;
 
PACKAGE BODY name IS
   -- Constructs implementation go here
   -- Function and procedure definitions go here
   ...

END name;
